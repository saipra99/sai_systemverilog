
class Packet;
Packet p;
